-- Library declarations
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;  -- Single library for arithmetic and conversion
use work.MyPackage.all;

-- Entity Declaration
entity fetchModule is
	port(
		hex0,hex1,hex2,hex3,hex4,hex5,hex6,hex7 	: out std_logic_vector(6 downto 0);
		leds 													: out std_logic_vector(3 downto 0);
		topclock,topreset 								: in std_logic
	
	); 
end fetchModule;

architecture bhv of fetchModule is

	
	-- TOP INSTRUCTION 
	-- TOP PC
	
	signal top_instruction , top_pcout : std_LOGIC_VECTOR(31 downto 0);

begin
	
	f1: fetch port map (
        PC_out             => top_pcout,
        instruction        => top_instruction,
        branch_addr        => X"00000000",
        jump_addr          => X"00000000",
        branch_decision    => '0', 				-- branch_des
        jump_decision      => '0',   			-- jump_des
        reset              => topreset,
        clock              => topclock
    );
	 leds <= top_pcout(3 downto 0);
	 
	 
u7: sevenSegement port map (
        bininput => top_instruction(31 downto 28),
        cathodes => hex7
    );
    u6: sevenSegement port map (
        bininput => top_instruction(27 downto 24),
        cathodes => hex6
    );
    u5: sevenSegement port map (
        bininput => top_instruction(23 downto 20),
        cathodes => hex5
    );
    u4: sevenSegement port map (
        bininput => top_instruction(19 downto 16),
        cathodes => hex4
    );
    u3: sevenSegement port map (
        bininput => top_instruction(15 downto 12),
        cathodes => hex3
    );
    u2: sevenSegement port map (
        bininput => top_instruction(11 downto 8),
        cathodes => hex2
    );
    u1: sevenSegement port map (
        bininput => top_instruction(7 downto 4),
        cathodes => hex1
    );
    u0: sevenSegement port map (
        bininput => top_instruction(3 downto 0),
        cathodes => hex0
    );
	
end bhv;