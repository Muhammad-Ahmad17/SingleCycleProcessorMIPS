library verilog;
use verilog.vl_types.all;
entity decodeModule_vlg_vec_tst is
end decodeModule_vlg_vec_tst;
